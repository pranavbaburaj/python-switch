module hello

pub fn hehe() {
	println("LOL")
}