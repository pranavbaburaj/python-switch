module std

// The std module that contains 
// a set of modules used for
// simple utilities
