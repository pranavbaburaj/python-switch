module std

// The std module 